module beers
import os

const (
  DB_USER = os.getenv('DB_USER')
  DB_PASS = os.getenv('DB_PASS')
  DB_NAME = os.getenv('DB_NAME')
  DB_HOST = os.getenv('DB_HOST')
  DB_PORT = os.getenv('DB_PORT')
)
